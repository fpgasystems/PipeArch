`ifndef GLM_COMMON
`define GLM_COMMON

// *************************************************************************
    //
    //   NUM_LOAD_CHANNELS
    //
    // *************************************************************************
    parameter NUM_LOAD_CHANNELS = 5;

    // *************************************************************************
    //
    //   NUM_WRITEBACK_CHANNELS
    //
    // *************************************************************************
    parameter NUM_WRITEBACK_CHANNELS = 2;

`endif // GLM_COMMON